library ieee;
use ieee.std_logic_1164.all;

package display7 is
    function segmentos7 (hex : std_logic_vector(3 downto 0))
                         return std_logic_vector;  -- 6 downto 0
end package;

package body display7 is
    function segmentos7 (hex : std_logic_vector(3 downto 0))
                         return std_logic_vector is
    begin
        case hex is
            when "0000" => return "1000000"; -- 0
            when "0001" => return "1111001"; -- 1
            when "0010" => return "0100100"; -- 2
            when "0011" => return "0110000"; -- 3
            when "0100" => return "0011001"; -- 4
            when "0101" => return "0010010"; -- 5
            when "0110" => return "0000010"; -- 6
            when "0111" => return "1111000"; -- 7
            when "1000" => return "0000000"; -- 8
            when "1001" => return "0010000"; -- 9
            when others => return "1111111"; -- tudo apagado
        end case;
    end;
end package body;
